module fa (input wire i0, i1, cin, output wire sum, cout);
   
endmodule

module addsub (input wire addsub, i0, i1, cin, output wire sumdiff, cout);
  
endmodule

module alu_slice (input wire [1:0] op, input wire i0, i1, cin, output wire o, cout);
  
endmodule

module alu (input wire [1:0] op, input wire [15:0] i0, i1,
    output wire [15:0] o, output wire cout);
  
endmodule
